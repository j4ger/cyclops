module cyclops_top;



endmodule

