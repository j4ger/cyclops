package interfaces;
  typedef struct {
    logic [7:0] red;
    logic [7:0] green;
    logic [7:0] blue;
    logic [7:0] depth;
  } pixel_t;



endpackage
